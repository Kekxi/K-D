// tf_ROM rom0(         
//                .clk(clk),
//                .A(tf_address),
//                .IREN(ren),
//                .KD_mode(KD_mode),

//                .Q(w));
module tf_ROM #(parameter addr_rom_width = 7,data_width = 36,depth_rom = 40)(  //addr_rom_width = 7---ROM 的地址宽度 2^7=128 Dilithium需要128个
    input clk,
    input [addr_rom_width-1:0] A,
    input IREN,
    input KD_mode,

    output reg [data_width-1:0] Q); 
    //需要区分k D 
    always@(posedge clk) begin
       if(IREN == 1'b1) begin
            if(KD_mode) begin
                case(A)
                    //Dilithium 256点24bit 去重后有128个24bit旋转因子  基2时 每轮蝶形运算需要1个24bit旋转因子 
                    //                                            十进制     二进制（23bit）           高11位（B） （D）  低12位（B） （D）
                    0:  Q <= 36'b00000000000000000000001; //W0:    1         00000000000000000000001   00000000000  0    000000000001 1   
                    1:  Q <= 36'b01010110110111010101111; //W1:    2846383   01010110110111010101111   01010110110  694  111010101111 3759  
                    2:  Q <= 36'b10111011001011000000011; //W2:    6133251   10111011001011000000011   10111011001  1481 011000000011 1539  
                    3:  Q <= 36'b00110110000001111001011; //W3:    1770443   00110110000001111001011   00110110000  432  001111001011 971  
                    4:  Q <= 36'b11001110100110111011111; //W4:    6770143   11001110100110111011111   11001110100  3300 110111011111 3583    
                    5:  Q <= 36'b01110010011001000100100; //W5:    3748388   01110010011001000100100   01110010011  1843 001000100100 548    
                    6:  Q <= 36'b11111000010111100001101; //W6:    8138509   11111000010111100001101   11111000010  4066 111100001101 3901    
                    7:  Q <= 36'b01011000000001010101110; //W7:    2884270   01011000000001010101110   01011000000  704  001010101110 686    
                    8:  Q <= 36'b00100001000101000010010; //W8:    1083922   00100001000101000010010   00100001000  264  101000010010 2578    
                    9:  Q <= 36'b10110100111111010111011; //W9:    5930683   10110100111111010111011   10110100111  1447 111010111011 3771    
                    10: Q <= 36'b01011010111111001001010; //W10:   2981450   01011010111111001001010   01011010111  727  111001001010 3626    
                    11: Q <= 36'b10110110110100001110001; //W11:   5990513   10110110110100001110001   10110110110  1462 100001110001 2145    
                    12: Q <= 36'b11001001111011111000100; //W12:   6617028   11001001111011111000100   11001001111  3215 011111000100 2020    
                    13: Q <= 36'b10110110000110010001100; //W13:   5966988   10110110000110010001100   10110110000  1456 110010001100 3116    
                    14: Q <= 36'b10110110100101000010111; //W14:   5982743   10110110100101000010111   10110110100  1460 101000010111 2607    
                    15: Q <= 36'b11100111100000001111010; //W15:   7585914   11100111100000001111010   11100111100  3676 000001111010 122    
                    16: Q <= 36'b10001011001011010000001; //W16:   4560513   10001011001011010000001   10001011001  2217 011010000001 1697    
                    17: Q <= 36'b01010000111111100110000; //W17:   2654000   01010000111111100110000   01010000111  647  111100110000 3920    
                    18: Q <= 36'b01100100001000111010011; //W18:   3281363   01100100001000111010011   01100100001  1601 000111010011 467    
                    19: Q <= 36'b01011010000011100111110; //W19:   2950974   01011010000011100111110   01011010000  720  011100111110 1854    
                    20: Q <= 36'b00110001101011001111100; //W20:   1627772   00110001101011001111100   00110001101  397  011001111100 1660    
                    21: Q <= 36'b00111011000100100011011; //W21:   1935643   00111011000100100011011   00111011000  472  100100011011 2379    
                    22: Q <= 36'b11100011101001111100110; //W22:   7459814   11100011101001111100110   11100011101  3629 001111100110 998    
                    23: Q <= 36'b11010000110001011100010; //W23:   6841058   11010000110001011100010   11010000110  3334 001011100010 722    
                    24: Q <= 36'b10100101011000000010101; //W24:   5419029   10100101011000000010101   10100101011  1323 000000010101 5    
                    25: Q <= 36'b00010000011111010001011; //W25:   540299    00010000011111010001011   00010000011  67   111010001011 3739    
                    26: Q <= 36'b10100110001001101001101; //W26:   5444429   10100110001001101001101   10100110001  1329 001101001101 861    
                    27: Q <= 36'b11111010001001111101110; //W27:   8197102   11111010001001111101110   11111010001  4001 001111101110 1022    
                    28: Q <= 36'b10111000101011010101111; //W28:   6051503   10111000101011010101111   10111000101  1477 011010101111 1711    
                    29: Q <= 36'b11110111010001111101101; //W29:   8102893   11110111010001111101101   11110111010  4026 001111101101 1021    
                    30: Q <= 36'b01000000001100000101110; //W30:   2103342   01000000001100000101110   01000000001  513  100000101110 2158    
                    31: Q <= 36'b00110001000001001011111; //W31:   1606239   00110001000001001011111   00110001000  392  001001011111 607    
                    32: Q <= 36'b10011001101000100111110; //W32:   5034302   10011001101000100111110   10011001101  2461 000100111110 318    
                    33: Q <= 36'b10100100001100111100011; //W33:   5380579   10100100001100111100011   10100100001  1313 100111100011 2531    
                    34: Q <= 36'b11011001011111101010001; //W34:   7126865   11011001011111101010001   11011001011  3531 111101010001 3937    
                    35: Q <= 36'b10100101000000001001101; //W35:   5406797   10100101000000001001101   10100101000  1320 000001001101 77    
                    36: Q <= 36'b01000100001111110111101; //W36:   2236349   01000100001111110111101   01000100001  545  111110111101 4061    
                    37: Q <= 36'b00010110001001011100100; //W37:   725732    00010110001001011100100   00010110001  89   001011100100 724    
                    38: Q <= 36'b11110000011000110011011; //W38:   7877019   11110000011000110011011   11110000011  3907 000110011011 411    
                    39: Q <= 36'b01110000010110010011001; //W39:   3681433   01110000010110010011001   01110000010  1794 110010011001 3209    
                    40: Q <= 36'b11111011101011100010101; //W40:   8247061   11111011101011100010101   11111011101  4061 011100010101 1813    
                    41: Q <= 36'b00010110010101000000001; //W41:   731649    00010110010101000000001   00010110010  90   101000000001 2561    
                    42: Q <= 36'b00100100010101110010100; //W42:   1190804   00100100010101110010100   00100100010  578  101110010100 2980    
                    43: Q <= 36'b11101010001110101111111; //W43:   7675263   11101010001110101111111   11101010001  3729 110101111111 3455    
                    44: Q <= 36'b01001001110001010001101; //W44:   2417293   01001001110001010001101   01001001110  590  001010001101 653    
                    45: Q <= 36'b10001111100001111111111; //W45:   4703231   10001111100001111111111   10001111100  2300 001111111111 1023    
                    46: Q <= 36'b01000100100000100101110; //W46:   2244910   01000100100000100101110   01000100100  548  000100101110 302    
                    47: Q <= 36'b11010110010101001000001; //W47:   7023169   11010110010101001000001   11010110010  3426 101001000001 1281     
                    48: Q <= 36'b10110110110001101011011; //W48:   5989211   10110110110001101011011   10110110110  1462 001101011011 859     
                    49: Q <= 36'b01100100110110011010100; //W49:   3304660   01100100110110011010100   01100100110  1606 110011010100 3252     
                    50: Q <= 36'b01000101111001111001001; //W50:   2290633   01000101111001111001001   01000101111  559  001111001001 969      
                    51: Q <= 36'b01101110110111110010000; //W51:   3633040   01101110110111110010000   01101110110  1774 111110010000 4000    
                    52: Q <= 36'b01011000101010101100110; //W52:   2905446   01011000101010101100110   01011000101  709  010101100110 1382    
                    53: Q <= 36'b00011110110000110100100; //W53:   1008036   00011110110000110100100   00011110110  246  000110100100 420    
                    54: Q <= 36'b10001000010000100010010; //W54:   4464914   10001000010000100010010   10001000010  2178 000100010010 274    
                    55: Q <= 36'b11111010110001110110101; //W55:   8217525   11111010110001110110101   11111010110  4022 001110110101 981    
                    56: Q <= 36'b10000111011011101111101; //W56:   4437885   10000111011011101111101   10000111011  2123 011101111101 1917    
                    57: Q <= 36'b11101100110011110111000; //W57:   7759800   11101100110011110111000   11101100110  3814 011110111000 2024    
                    58: Q <= 36'b01100101001010100010000; //W58:   3314960   01100101001010100010000   01100101001  1609 010100010000 1344    
                    59: Q <= 36'b10110110111011101010000; //W59:   5994320   10110110111011101010000   10110110111  1463 011101010000 1872    
                    60: Q <= 36'b10000001111110010100101; //W60:   4258981   10000001111110010100101   10000001111  2063 110010100101 3237    
                    61: Q <= 36'b10001100101110100101100; //W61:   4611372   10001100101110100101100   10001100101  2245 110100101100 3436    
                    62: Q <= 36'b10011010010110110000010; //W62:   5057922   10011010010110110000010   10011010010  2474 110110000010 3458    
                    63: Q <= 36'b11100111010000101111111; //W63:   7577983   11100111010000101111111   11100111010  3674 000101111111 383    
                    64: Q <= 36'b10001111101011110001000; //W64:   4708232   10001111101011110001000   10001111101  2301 011110001000 1992     
                    65: Q <= 36'b11001111110000001101001; //W65:   6807657   11001111110000001101001   11001111110  3326 000001101001 105     
                    66: Q <= 36'b11101010011010101011010; //W66:   7681370   11101010011010101011010   11101010011  3731 010101011010 1386     
                    67: Q <= 36'b10101111011010101010011; //W67:   5748051   10101111011010101010011   10101111011  1403 010101010011 1363    
                    68: Q <= 36'b10100101010000101011100; //W68:   5415260   10100101010000101011100   10100101010  1322 000101011100 348    
                    69: Q <= 36'b01010101101111100010011; //W69:   2809619   01010101101111100010011   01010101101  685  111100010011 3891    
                    70: Q <= 36'b00101001011001100010111; //W70:   1356567   00101001011001100010111   00101001011  683  001100010111 775     
                    71: Q <= 36'b10011100111100010100100; //W71:   5142692   10011100111100010100100   10011100111  2535 100010100100 2212     
                    72: Q <= 36'b11001010101101000100000; //W72:   6642208   11001010101101000100000   11001010101  3237 101000100000 2624     
                    73: Q <= 36'b01001010101110111101101; //W73:   2448877   01001010101110111101101   01001010101  597  110111101101 3573     
                    74: Q <= 36'b00000110110111011011000; //W74:   224984    00000110110111011011000   00000110110  54   111011011000 3816     
                    75: Q <= 36'b11011010010101000001000; //W75:   7154184   11011010010101000001000   11011010010  3538 101000001000 2568     
                    76: Q <= 36'b01011110000010100100001; //W76:   3081505   01011110000010100100001   01011110000  752  010100100001 1313     
                    77: Q <= 36'b01110001111011111010100; //W77:   3733460   01110001111011111010100   01110001111  1855 011111010100 2004     
                    78: Q <= 36'b11101010100101111101101; //W78:   7687149   11101010100101111101101   11101010100  3732 101111101101 3037     
                    79: Q <= 36'b01101001011011100000101; //W79:   3454725   01101001011011100000101   01101001011  1683 011100000101 1797     
                    80: Q <= 36'b10010000010001101000100; //W80:   4727620   10010000010001101000100   10010000010  2306 001101000100 836    
                    81: Q <= 36'b10110001011001100001101; //W81:   5813005   10110001011001100001101   10110001011  1427 001100001101 781    
                    82: Q <= 36'b01010101100100111110100; //W82:   2804212   01010101100100111110100   01010101100  684  100111110100 2548    
                    83: Q <= 36'b11101011101001001001001; //W83:   7721545   11101011101001001001001   11101011101  3773 001001001001 585    
                    84: Q <= 36'b11000110000000110111111; //W84:   6488511   11000110000000110111111   11000110000  3168 000110111111 447    
                    85: Q <= 36'b10011111111011101100001; //W85:   5240673   10011111111011101100001   10011111111  2559 011101100001 1889    
                    86: Q <= 36'b00000010101000000110110; //W86:   86070     00000010101000000110110   00000010101  21   000000110110 54    
                    87: Q <= 36'b10100101010110101110011; //W87:   5418355   10100101010110101110011   10100101010  1322 110101110011 3443    
                    88: Q <= 36'b00100101011011101011010; //W88:   1226586   00100101011011101011010   00100101011  587  011101011010 1898    
                    89: Q <= 36'b01000100011000111110101; //W89:   2241013   01000100011000111110101   01000100011  547  000111110101 501    
                    90: Q <= 36'b10010000110101011000111; //W90:   4745927   10010000110101011000111   10010000110  2302 101011000111 2767    
                    91: Q <= 36'b01110110010001010110010; //W91:   3875506   01110110010001010110010   01110110010  1890 001010110010 690    
                    92: Q <= 36'b10100100100010011010101; //W92:   5391573   10100100100010011010101   10100100100  1316 010011010101 1237    
                    93: Q <= 36'b10000010110100010100110; //W93:   4286630   10000010110100010100110   10000010110  2150 100010100110 2214    
                    94: Q <= 36'b10110100101010111100010; //W94:   5920226   10110100101010111100010   10110100101  1445 010111100010 754    
                    95: Q <= 36'b00111011010110011100000; //W95:   1944800   00111011010110011100000   00111011010  474  110011100000 3296    
                    96: Q <= 36'b00000011011001110101001; //W96:   111529    00000011011001110101001   00000011011  27   001110101001 937    
                    97: Q <= 36'b11001001100010110110100; //W97:   6604212   11001001100010110110100   11001001100  3180 010110110100 1460    
                    98: Q <= 36'b00110001000010111100111; //W98:   1607143   00110001000010111100111   00110001000  392  010111100111 759    
                    99: Q <= 36'b11110001010001011010110; //W99:   7906006   11110001010001011010110   11110001010  3898 001011010110 726    
                    100:Q <= 36'b11000000011000111110111; //W100： 6304247   11000000011000111110111   11000000011  3075 000111110111 503   
                    101:Q <= 36'b01110000111100111100111; //W101： 3701223   01110000111100111100111   01110000111  1799 100111100111 2551   
                    102:Q <= 36'b01010010000000101110111; //W102： 2687351   01010010000000101110111   01010010000  656  000101110111 375   
                    103:Q <= 36'b11000111100000111010110; //W103： 6537686   11000111100000111010110   11000111100  3196 000111010110 470   
                    104:Q <= 36'b00101110101111000110111; //W104： 1531447   00101110101111000110111   00101110101  757  111000110111 3647    
                    105:Q <= 36'b00100011010111100111001; //W105： 1158969   00100011010111100111001   00100011010  570  111100111001 3993    
                    106:Q <= 36'b11111101101001001111001; //W106： 8311417   11111101101001001111001   11111101101  4061 001001111001 633    
                    107:Q <= 36'b01111011001011100001011; //W107： 4036363   01111011001011100001011   01111011001  1977 011100001011 1803    
                    108:Q <= 36'b01001011001100100010010; //W108： 2464018   01001011001100100010010   01001011001  601  100100010010 2338    
                    109:Q <= 36'b01010010111000110010111; //W109： 2716055   01010010111000110010111   01010010111  663  000110010111 407    
                    110:Q <= 36'b01110000010111010010010; //W110： 3681938   01110000010111010010010   01110000010  1794 111010010010 3730    
                    111:Q <= 36'b00010101111001010111000; //W111： 717496    00010101111001010111000   00010101111  95   001010111000 696    
                    112:Q <= 36'b01100011101000101001000; //W112： 3264840   01100011101000101001000   01100011101  1581 000101001000 328    
                    113:Q <= 36'b10101000110001111000000; //W113： 5530560   10101000110001111000000   10101000110  1350 001111000000 992    
                    114:Q <= 36'b01000010110110111101011; //W114： 2190827   01000010110110111101011   01000010110  534  110111101011 3563    
                    115:Q <= 36'b01011110001000100011101; //W115： 3084573   01011110001000100011101   01011110001  753  000100011101 285    
                    116:Q <= 36'b11111110010001110101010; //W116： 8332202   11111110010001110101010   11111110010  4066 001110101010 954    
                    117:Q <= 36'b01110111111110110111110; //W117： 3931582   01110111111110110111110   01110111111  1919 110110111110 3518    
                    118:Q <= 36'b10101110110101101100111; //W118： 5729127   10101110110101101100111   10101110110  1398 101101100111 2927    
                    119:Q <= 36'b01000111110101111100101; //W119： 2354149   01000111110101111100101   01000111110  574  101111100101 3045    
                    120:Q <= 36'b01000011011001010010000; //W120： 2208400   01000011011001010010000   01000011011  523  001010010000 656    
                    121:Q <= 36'b11100101100100000110001; //W121： 7522353   11100101100100000110001   11100101100  3660 100000110001 2145    
                    122:Q <= 36'b01100011100000000000001; //W122： 3260417   01100011100000000000001   01100011100  1580 000000000001 1    
                    123:Q <= 36'b10110001110101011101101; //W123： 5827309   10110001110101011101101   10110001110  1422 101011101101 2781    
                    124:Q <= 36'b01101011111100111111001; //W124： 3537401   01101011111100111111001   01101011111  1727 100111111001 2553   
                    125:Q <= 36'b10011000001011101100110; //W125： 4986726   10011000001011101100110   10011000001  2433 011101100110 1894   
                    126:Q <= 36'b01010110111000010000110; //W126： 2846854   01010110111000010000110   01010110111  695  000010000110 134   
                    127:Q <= 36'b00001000000011110011100; //W127： 264092    00001000000011110011100   00001000000  64   011110011100 1956 
                endcase   
            end else begin //Kyber
                case(A) 
                  //                                                        w1     w2   w3
                  0:  Q <= 36'b010010010010100000111110010100001111;   //   1170  2110 1295        010010010010   100000111110   010100001111
                  1:  Q <= 36'b010000100100011000011000011110111100;   //   1060  1560 1980        010000100100   011000011000   011110111100
                  2:  Q <= 36'b010110101001010010110011011101111100;   //   1449  1203 1916        010110101001   010010110011   011101111100
                  3:  Q <= 36'b011011101111000000111001000110100011;   //   1775    57  419        011011101111   000000111001   000110100011
                  4:  Q <= 36'b100000010100010001101101000000110001;   //   2068  1133   49        100000010100   010001101101   000000110001
                  5:  Q <= 36'b010110001110001010011011011101101010;   //   1422   667 1898        010110001110   001010011011   011101101010
                  6:  Q <= 36'b100001011101000100000100000110000011;   //   2141   260  387        100001011101   000100000100   000110000011
                  7:  Q <= 36'b100010000110100010111100001001010000;   //   2182  2236  592        100010000110   100010111100   001001010000
                  8:  Q <= 36'b010100111101100000100000000001000010;   //   1341  2080   66        010100111101   100000100000   000001000010
                  9:  Q <= 36'b000110000111011010010001010011000111;   //    391  1681 1223        000110000111   011010010001   010011000111
                  10: Q <= 36'b011100011001010101111010001010110110;   //   1817  1402  694        011100011001   010101111010   001010110110
                  11: Q <= 36'b000110010010011110101001010010101101;   //    402  1961 1197        000110010010   011110101001   010010101101
                  12: Q <= 36'b010100001111010001000111000101100110;   //   1295  1095  358        010100001111   010001000111   000101100110
                  13: Q <= 36'b011110111100010011001110100001000011;   //   1980  1230 2115        011110111100   010011001110   100001000011
                  14: Q <= 36'b011101111100010010111100000000111101;   //   1916  1212   61        011101111100   010010111100   000000111101
                  15: Q <= 36'b000110100011001010011000000000010010;   //    419   664   18        000110100011   001010011000   000000010010
                  16: Q <= 36'b000000110001100010110000100000010110;   //     49  2224 2070        000000110001   100010110000   100000010110
                  17: Q <= 36'b011101101010000000000110001011110101;   //   1898     6  757        011101101010   000000000110   001011110101
                  18: Q <= 36'b000110000011010111000101001010011100;   //    387  1477  668        000110000011   010111000101   001010011100
                  19: Q <= 36'b001001010000001111000101001011001000;   //    592   965  712        001001010000   001111000101   001011001000
                  20: Q <= 36'b010011010100010010010010100000111110;   //   1236  1170  2110       010011010100   010010010010   100000111110
                  21: Q <= 36'b010010011010010000100100011000011000;   //   1178  1060  1560       010010011010   010000100100   011000011000
                  22: Q <= 36'b000100101100010110101001010010110011;   //    300  1449  1203       000100101100   010110101001   010010110011
                  23: Q <= 36'b000110111101011011101111000000111001;   //    445  1775    57       000110111101   011011101111   000000111001
                  24: Q <= 36'b000110010111100000010100010001101101;   //    407  2068  1133       000110010111   100000010100   010001101101
                  25: Q <= 36'b010011100001010110001110001010011011;   //   1249  1422   667       010011100001   010110001110   001010011011
                  26: Q <= 36'b100000011010100001011101000100000100;   //   2074  2141   260       100000011010   100001011101   000100000100
                  27: Q <= 36'b000111010001100010000110100010111100;   //    465  2182  2236       000111010001   100010000110   100010111100
                  28: Q <= 36'b010011000001010100111101100000100000;   //   1217  1341  2080       010011000001   010100111101   100000100000
                  29: Q <= 36'b000101010010000110000111011010010001;   //    338   391  1681       000101010010   000110000111   011010010001
                  30: Q <= 36'b010010101001011100011001010101111010;   //   1193  1817  1402       010010101001   011100011001   010101111010
                  31: Q <= 36'b001101110111000110010010011110101001;   //    887   402  1961       001101110111   000110010010   011110101001
                  32: Q <= 36'b100000111110010100001111010001000111;   //   2110  1295  1095       100000111110   010100001111   010001000111
                  33: Q <= 36'b011000011000011110111100010011001110;   //   1560  1980  1230       011000011000   011110111100   010011001110
                  34: Q <= 36'b010010110011011101111100010010111100;   //   1203  1916  1212       010010110011   011101111100   010010111100
                  35: Q <= 36'b000000111001000110100011001010011000;   //     57   419   664       000000111001   000110100011   001010011000
                  36: Q <= 36'b010001101101000000110001100010110000;   //   1133    49  2224       010001101101   000000110001   100010110000
                  37: Q <= 36'b001010011011011101101010000000000110;   //    667  1898     6       001010011011   011101101010   000000000110
                  38: Q <= 36'b000100000100000110000011010111000101;   //    260   387  1477       000100000100   000110000011   010111000101
                  39: Q <= 36'b100010111100001001010000001111000101;   //   2236   592   965       100010111100   001001010000   001111000101
                  40: Q <= 36'b100000100000000001000010010110101001;   //   2080    66  1449       100000100000   000001000010   010110101001
                  41: Q <= 36'b011010010001010011000111011011101111;   //   1681  1223  1775       011010010001   010011000111   011011101111

                    // //如果按照这种方式 旋转因子取的时候需要映射 因为点数相对较少 可以不复用旋转因子 1个地址中存基4蝶形运算的3个旋转因子
                    // //Kyber 128点 12bit 先算1个基2阶段 旋转因子1个（W0） 再算3个基4阶段 基4时蝶形运算需要3个旋转因子，2个重复  实际存2个 重复取即可 （但ROM位宽36 也会浪费12）
                    // //                                                   十进制           二进制（12bit）
                    // 0:  Q <= 36'b100000111110010100001111;   //W1  W0 :   2110 1295        100000111110   010100001111
                    // 1:  Q <= 36'b011000011000011110111100;   //W3  W2 :   1560 1980        011000011000   011110111100
                    // 2:  Q <= 36'b010010110011011101111100;   //W5  W4 :   1203 1916        010010110011   011101111100
                    // 3:  Q <= 36'b000000111001000110100011;   //W7  W6 :     57  419        000000111001   000110100011
                    // 4:  Q <= 36'b010001101101000000110001;   //W9  W8 :   1133   49        010001101101   000000110001
                    // 5:  Q <= 36'b001010011011011101101010;   //W11 W10:    667 1898        001010011011   011101101010
                    // 6:  Q <= 36'b000100000100000110000011;   //W13 W12:    260  387        000100000100   000110000011
                    // 7:  Q <= 36'b100010111100001001010000;   //W15 W14:   2236  592        100010111100   001001010000
                    // 8:  Q <= 36'b100000100000000001000010;   //W17 W16:   2080   66        100000100000   000001000010
                    // 9:  Q <= 36'b011010010001010011000111;   //W19 W18    1681 1223        011010010001   010011000111
                    // 10: Q <= 36'b010101111010001010110110;   //W21 W20:   1402  694        010101111010   001010110110
                    // 11: Q <= 36'b011110101001010010101101;   //W23 W22:   1961 1197        011110101001   010010101101
                    // 12: Q <= 36'b010001000111000101100110;   //W25 W24:   1095  358        010001000111   000101100110
                    // 13: Q <= 36'b010011001110100001000011;   //W27 W26:   1230 2115        010011001110   100001000011
                    // 14: Q <= 36'b010010111100000000111101;   //W29 W28:   1212   61        010010111100   000000111101
                    // 15: Q <= 36'b001010011000000000010010;   //W31 W30:    664   18        001010011000   000000010010
                    // 16: Q <= 36'b100010110000100000010110;   //W33 W32:   2224 2070        100010110000   100000010110
                    // 17: Q <= 36'b000000000110001011110101;   //W35 W34:      6  757        000000000110   001011110101
                    // 18: Q <= 36'b010111000101001010011100;   //W37 W36:   1477  668        010111000101   001010011100
                    // 19: Q <= 36'b001111000101001011001000;   //W39 W38:    965  712        001111000101   001011001000
                    // 20: Q <= 36'b010011010100010010010010;   //W41 W40:   1236 1170        010011010100   010010010010
                    // 21: Q <= 36'b010010011010010000100100;   //W43 W42:   1178 1060        010010011010   010000100100
                    // 22: Q <= 36'b000100101100010110101001;   //W45 W44:    300 1449        000100101100   010110101001
                    // 23: Q <= 36'b000110111101011011101111;   //W47 W46:    445 1775        000110111101   011011101111
                    // 24: Q <= 36'b000110010111100000010100;   //W49 W48:    407 2068        000110010111   100000010100
                    // 25: Q <= 36'b010011100001010110001110;   //W51 W50:   1249 1422        010011100001   010110001110
                    // 26: Q <= 36'b100000011010100001011101;   //W53 W52:   2074 2141        100000011010   100001011101
                    // 27: Q <= 36'b000111010001100010000110;   //W55 W54:    465 2182        000111010001   100010000110
                    // 28: Q <= 36'b010011000001010100111101;   //W57 W56:   1217 1341        010011000001   010100111101
                    // 29: Q <= 36'b000101010010000110000111;   //W59 W58:    338  391        000101010010   000110000111
                    // 30: Q <= 36'b010010101001011100011001;   //W61 W60:   1193 1817        010010101001   011100011001
                    // 31: Q <= 36'b001101110111000110010010;   //W63 W62:    887  402        001101110111   000110010010

                endcase
            end
        end         
    end
endmodule